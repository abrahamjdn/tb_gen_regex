    
    
    module test  (
        input a,b,c,d,
    input [     0         :  31] ye, f,
    input sal_0,
    output sal_1,
    output [3:0] sal_2, // otro ejemplo
    //salidas de todo
/* comentario */ output k,
/*comentario extra*/

input zz,yy,ss,dd,
/*
    comentario de varias 
    lineas
*/ output test123456,
/*
pruebas
*/
/*
mas pruebas
*/
    output [3:0 ] sal_3,

    output [ 3 : 0 ] sal_4,sal_5,        sal_6,
    input clk       
    );
    /*
    Bla Bla Bla
    Bla Bla Bla
    */
endmodule